module not_gate (
    input wire a,
    output wire b
);

    assign b = ~a;

endmodule